module binbcd (

	input logic [7:0] bin,
	output logic [3:0] bcd0,
	output logic [3:0] bcd1);
	
	always @(*)
		case(bin)
		
			8'b00000000: begin
					  bcd1 = 4'b0000;
					  bcd0 = 4'b0000;
					  end

			8'b00000001: begin
					  bcd1 = 4'b0000;
					  bcd0 = 4'b0001;
					  end

			8'b00000010: begin
					  bcd1 = 4'b0000;
					  bcd0 = 4'b0010;
					  end

			8'b00000011: begin
					  bcd1 = 4'b0000;
					  bcd0 = 4'b0011;
					  end

			8'b00000100: begin
					  bcd1 = 4'b0000;
					  bcd0 = 4'b0100;
					  end

			8'b00000101: begin
					  bcd1 = 4'b0000;
					  bcd0 = 4'b0101;
					  end

			8'b00000110: begin
					  bcd1 = 4'b0000;
					  bcd0 = 4'b0110;
					  end

			8'b00000111: begin
					  bcd1 = 4'b0000;
					  bcd0 = 4'b0111;
					  end

			8'b00001000: begin
					  bcd1 = 4'b0000;
					  bcd0 = 4'b1000;
					  end

			8'b00001001: begin
					  bcd1 = 4'b0000;
					  bcd0 = 4'b1001;
					  end

			8'b00001010: begin
					  bcd1 = 4'b0001;
					  bcd0 = 4'b0000;
					  end

			8'b00001011: begin
					  bcd1 = 4'b0001;
					  bcd0 = 4'b0001;
					  end

			8'b00001100: begin
					  bcd1 = 4'b0001;
					  bcd0 = 4'b0010;
					  end

			8'b00001101: begin
					  bcd1 = 4'b0001;
					  bcd0 = 4'b0011;
					  end

			8'b00001110: begin
					  bcd1 = 4'b0001;
					  bcd0 = 4'b0100;
					  end

			8'b00001111: begin
					  bcd1 = 4'b0001;
					  bcd0 = 4'b0101;
					  end

			8'b00010000: begin
					  bcd1 = 4'b0001;
					  bcd0 = 4'b0110;
					  end

			8'b00010001: begin
					  bcd1 = 4'b0001;
					  bcd0 = 4'b0111;
					  end

			8'b00010010: begin
					  bcd1 = 4'b0001;
					  bcd0 = 4'b1000;
					  end

			8'b00010011: begin
					  bcd1 = 4'b0001;
					  bcd0 = 4'b1001;
					  end

			8'b00010100: begin
					  bcd1 = 4'b0010;
					  bcd0 = 4'b0000;
					  end

			8'b00010101: begin
					  bcd1 = 4'b0010;
					  bcd0 = 4'b0001;
					  end

			8'b00010110: begin
					  bcd1 = 4'b0010;
					  bcd0 = 4'b0010;
					  end

			8'b00010111: begin
					  bcd1 = 4'b0010;
					  bcd0 = 4'b0011;
					  end

			8'b00011000: begin
					  bcd1 = 4'b0010;
					  bcd0 = 4'b0100;
					  end

			8'b00011001: begin
					  bcd1 = 4'b0010;
					  bcd0 = 4'b0101;
					  end

			8'b00011010: begin
					  bcd1 = 4'b0010;
					  bcd0 = 4'b0110;
					  end

			8'b00011011: begin
					  bcd1 = 4'b0010;
					  bcd0 = 4'b0111;
					  end

			8'b00011100: begin
					  bcd1 = 4'b0010;
					  bcd0 = 4'b1000;
					  end

			8'b00011101: begin
					  bcd1 = 4'b0010;
					  bcd0 = 4'b1001;
					  end

			8'b00011110: begin
					  bcd1 = 4'b0011;
					  bcd0 = 4'b0000;
					  end

			8'b00011111: begin
					  bcd1 = 4'b0011;
					  bcd0 = 4'b0001;
					  end

			8'b00100000: begin
					  bcd1 = 4'b0011;
					  bcd0 = 4'b0010;
					  end

			8'b00100001: begin
					  bcd1 = 4'b0011;
					  bcd0 = 4'b0011;
					  end

			8'b00100010: begin
					  bcd1 = 4'b0011;
					  bcd0 = 4'b0100;
					  end

			8'b00100011: begin
					  bcd1 = 4'b0011;
					  bcd0 = 4'b0101;
					  end

			8'b00100100: begin
					  bcd1 = 4'b0011;
					  bcd0 = 4'b0110;
					  end

			8'b00100101: begin
					  bcd1 = 4'b0011;
					  bcd0 = 4'b0111;
					  end

			8'b00100110: begin
					  bcd1 = 4'b0011;
					  bcd0 = 4'b1000;
					  end

			8'b00100111: begin
					  bcd1 = 4'b0011;
					  bcd0 = 4'b1001;
					  end

			8'b00101000: begin
					  bcd1 = 4'b0100;
					  bcd0 = 4'b0000;
					  end

			8'b00101001: begin
					  bcd1 = 4'b0100;
					  bcd0 = 4'b0001;
					  end

			8'b00101010: begin
					  bcd1 = 4'b0100;
					  bcd0 = 4'b0010;
					  end

			8'b00101011: begin
					  bcd1 = 4'b0100;
					  bcd0 = 4'b0011;
					  end

			8'b00101100: begin
					  bcd1 = 4'b0100;
					  bcd0 = 4'b0100;
					  end

			8'b00101101: begin
					  bcd1 = 4'b0100;
					  bcd0 = 4'b0101;
					  end

			8'b00101110: begin
					  bcd1 = 4'b0100;
					  bcd0 = 4'b0110;
					  end

			8'b00101111: begin
					  bcd1 = 4'b0100;
					  bcd0 = 4'b0111;
					  end

			8'b00110000: begin
					  bcd1 = 4'b0100;
					  bcd0 = 4'b1000;
					  end

			8'b00110001: begin
					  bcd1 = 4'b0100;
					  bcd0 = 4'b1001;
					  end

			8'b00110010: begin
					  bcd1 = 4'b0101;
					  bcd0 = 4'b0000;
					  end

			8'b00110011: begin
					  bcd1 = 4'b0101;
					  bcd0 = 4'b0001;
					  end

			8'b00110100: begin
					  bcd1 = 4'b0101;
					  bcd0 = 4'b0010;
					  end

			8'b00110101: begin
					  bcd1 = 4'b0101;
					  bcd0 = 4'b0011;
					  end

			8'b00110110: begin
					  bcd1 = 4'b0101;
					  bcd0 = 4'b0100;
					  end

			8'b00110111: begin
					  bcd1 = 4'b0101;
					  bcd0 = 4'b0101;
					  end

			8'b00111000: begin
					  bcd1 = 4'b0101;
					  bcd0 = 4'b0110;
					  end

			8'b00111001: begin
					  bcd1 = 4'b0101;
					  bcd0 = 4'b0111;
					  end

			8'b00111010: begin
					  bcd1 = 4'b0101;
					  bcd0 = 4'b1000;
					  end

			8'b00111011: begin
					  bcd1 = 4'b0101;
					  bcd0 = 4'b1001;
					  end

			8'b00111100: begin
					  bcd1 = 4'b0110;
					  bcd0 = 4'b0000;
					  end

			8'b00111101: begin
					  bcd1 = 4'b0110;
					  bcd0 = 4'b0001;
					  end

			8'b00111110: begin
					  bcd1 = 4'b0110;
					  bcd0 = 4'b0010;
					  end

			8'b00111111: begin
					  bcd1 = 4'b0110;
					  bcd0 = 4'b0011;
					  end

			8'b01000000: begin
					  bcd1 = 4'b0110;
					  bcd0 = 4'b0100;
					  end

			8'b01000001: begin
					  bcd1 = 4'b0110;
					  bcd0 = 4'b0101;
					  end

			8'b01000010: begin
					  bcd1 = 4'b0110;
					  bcd0 = 4'b0110;
					  end

			8'b01000011: begin
					  bcd1 = 4'b0110;
					  bcd0 = 4'b0111;
					  end

			8'b01000100: begin
					  bcd1 = 4'b0110;
					  bcd0 = 4'b1000;
					  end

			8'b01000101: begin
					  bcd1 = 4'b0110;
					  bcd0 = 4'b1001;
					  end

			8'b01000110: begin
					  bcd1 = 4'b0111;
					  bcd0 = 4'b0000;
					  end

			8'b01000111: begin
					  bcd1 = 4'b0111;
					  bcd0 = 4'b0001;
					  end

			8'b01001000: begin
					  bcd1 = 4'b0111;
					  bcd0 = 4'b0010;
					  end

			8'b01001001: begin
					  bcd1 = 4'b0111;
					  bcd0 = 4'b0011;
					  end

			8'b01001010: begin
					  bcd1 = 4'b0111;
					  bcd0 = 4'b0100;
					  end

			8'b01001011: begin
					  bcd1 = 4'b0111;
					  bcd0 = 4'b0101;
					  end

			8'b01001100: begin
					  bcd1 = 4'b0111;
					  bcd0 = 4'b0110;
					  end

			8'b01001101: begin
					  bcd1 = 4'b0111;
					  bcd0 = 4'b0111;
					  end

			8'b01001110: begin
					  bcd1 = 4'b0111;
					  bcd0 = 4'b1000;
					  end

			8'b01001111: begin
					  bcd1 = 4'b0111;
					  bcd0 = 4'b1001;
					  end

			8'b01010000: begin
					  bcd1 = 4'b1000;
					  bcd0 = 4'b0000;
					  end

			8'b01010001: begin
					  bcd1 = 4'b1000;
					  bcd0 = 4'b0001;
					  end

			8'b01010010: begin
					  bcd1 = 4'b1000;
					  bcd0 = 4'b0010;
					  end

			8'b01010011: begin
					  bcd1 = 4'b1000;
					  bcd0 = 4'b0011;
					  end

			8'b01010100: begin
					  bcd1 = 4'b1000;
					  bcd0 = 4'b0100;
					  end

			8'b01010101: begin
					  bcd1 = 4'b1000;
					  bcd0 = 4'b0101;
					  end

			8'b01010110: begin
					  bcd1 = 4'b1000;
					  bcd0 = 4'b0110;
					  end

			8'b01010111: begin
					  bcd1 = 4'b1000;
					  bcd0 = 4'b0111;
					  end

			8'b01011000: begin
					  bcd1 = 4'b1000;
					  bcd0 = 4'b1000;
					  end

			8'b01011001: begin
					  bcd1 = 4'b1000;
					  bcd0 = 4'b1001;
					  end

			8'b01011010: begin
					  bcd1 = 4'b1001;
					  bcd0 = 4'b0000;
					  end

			8'b01011011: begin
					  bcd1 = 4'b1001;
					  bcd0 = 4'b0001;
					  end

			8'b01011100: begin
					  bcd1 = 4'b1001;
					  bcd0 = 4'b0010;
					  end

			8'b01011101: begin
					  bcd1 = 4'b1001;
					  bcd0 = 4'b0011;
					  end

			8'b01011110: begin
					  bcd1 = 4'b1001;
					  bcd0 = 4'b0100;
					  end

			8'b01011111: begin
					  bcd1 = 4'b1001;
					  bcd0 = 4'b0101;
					  end

			8'b01100000: begin
					  bcd1 = 4'b1001;
					  bcd0 = 4'b0110;
					  end

			8'b01100001: begin
					  bcd1 = 4'b1001;
					  bcd0 = 4'b0111;
					  end

			8'b01100010: begin
					  bcd1 = 4'b1001;
					  bcd0 = 4'b1000;
					  end

			8'b01100011: begin
					  bcd1 = 4'b1001;
					  bcd0 = 4'b1001;
					  end
		endcase

endmodule